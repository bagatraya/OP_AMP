magic
tech sky130A
magscale 1 2
timestamp 1729197635
<< nwell >>
rect 324 -1596 1124 912
<< nsubdiff >>
rect 360 842 420 876
rect 1028 842 1088 876
rect 360 816 394 842
rect 1054 816 1088 842
rect 360 -1526 394 -1500
rect 1054 -1526 1088 -1500
rect 360 -1560 420 -1526
rect 1028 -1560 1088 -1526
<< nsubdiffcont >>
rect 420 842 1028 876
rect 360 -1500 394 816
rect 1054 -1500 1088 816
rect 420 -1560 1028 -1526
<< poly >>
rect 508 259 538 289
rect 447 243 538 259
rect 447 209 463 243
rect 497 209 538 243
rect 447 193 538 209
rect 912 259 942 301
rect 912 243 1004 259
rect 912 209 954 243
rect 988 209 1004 243
rect 912 193 1004 209
rect 508 -233 538 -203
rect 445 -249 538 -233
rect 445 -283 461 -249
rect 495 -283 538 -249
rect 445 -299 538 -283
rect 912 -234 942 -202
rect 912 -250 1004 -234
rect 912 -284 954 -250
rect 988 -284 1004 -250
rect 596 -397 696 -299
rect 754 -397 854 -299
rect 912 -300 1004 -284
rect 446 -413 538 -397
rect 446 -447 462 -413
rect 496 -447 538 -413
rect 446 -463 538 -447
rect 508 -494 538 -463
rect 912 -413 1003 -397
rect 912 -447 953 -413
rect 987 -447 1003 -413
rect 912 -463 1003 -447
rect 912 -494 942 -463
rect 446 -906 538 -890
rect 446 -940 462 -906
rect 496 -940 538 -906
rect 446 -956 538 -940
rect 508 -987 538 -956
rect 912 -906 1004 -890
rect 912 -940 954 -906
rect 988 -940 1004 -906
rect 912 -956 1004 -940
rect 912 -987 942 -956
<< polycont >>
rect 463 209 497 243
rect 954 209 988 243
rect 461 -283 495 -249
rect 954 -284 988 -250
rect 462 -447 496 -413
rect 953 -447 987 -413
rect 462 -940 496 -906
rect 954 -940 988 -906
<< locali >>
rect 360 842 420 876
rect 1028 842 1088 876
rect 360 816 394 842
rect 1054 816 1088 842
rect 462 243 497 302
rect 954 243 988 302
rect 447 209 463 243
rect 497 209 513 243
rect 938 209 954 243
rect 988 209 1004 243
rect 461 -249 495 -190
rect 445 -283 461 -249
rect 495 -283 511 -249
rect 954 -250 988 -190
rect 938 -284 954 -250
rect 988 -284 1004 -250
rect 446 -447 462 -413
rect 496 -447 512 -413
rect 937 -447 953 -413
rect 987 -447 1003 -413
rect 462 -506 496 -447
rect 954 -506 989 -447
rect 446 -940 462 -906
rect 496 -940 512 -906
rect 938 -940 954 -906
rect 988 -940 1004 -906
rect 462 -999 496 -940
rect 954 -999 988 -940
rect 360 -1526 394 -1500
rect 1054 -1526 1088 -1500
rect 360 -1560 420 -1526
rect 1028 -1560 1088 -1526
<< viali >>
rect 557 876 767 877
rect 557 842 767 876
rect 463 209 497 243
rect 954 209 988 243
rect 461 -283 495 -249
rect 954 -284 988 -250
rect 462 -447 496 -413
rect 953 -447 987 -413
rect 462 -940 496 -906
rect 954 -940 988 -906
<< metal1 >>
rect 545 877 779 883
rect 545 842 557 877
rect 767 842 779 877
rect 545 836 779 842
rect 496 804 1002 808
rect 496 748 941 804
rect 997 748 1007 804
rect 496 418 556 748
rect 860 478 994 490
rect 456 289 590 418
rect 687 302 697 478
rect 753 302 763 478
rect 860 302 901 478
rect 953 302 994 478
rect 860 290 994 302
rect 462 249 497 289
rect 451 243 509 249
rect 451 209 463 243
rect 497 209 509 243
rect 451 203 509 209
rect 620 171 672 243
rect 760 200 770 252
rect 838 200 848 252
rect 954 249 988 290
rect 942 243 1000 249
rect 942 209 954 243
rect 988 209 1000 243
rect 942 203 1000 209
rect 620 119 830 171
rect 602 36 612 88
rect 680 36 690 88
rect 778 57 830 119
rect 456 -14 590 -2
rect 860 -14 994 -2
rect 443 -190 453 -14
rect 505 -190 590 -14
rect 687 -190 697 -14
rect 753 -190 763 -14
rect 860 -190 943 -14
rect 999 -190 1009 -14
rect 456 -202 590 -190
rect 860 -202 994 -190
rect 461 -243 495 -202
rect 449 -249 507 -243
rect 954 -244 988 -202
rect 449 -283 461 -249
rect 495 -283 507 -249
rect 449 -289 507 -283
rect 942 -250 1000 -244
rect 942 -284 954 -250
rect 988 -284 1000 -250
rect 942 -290 1000 -284
rect 450 -413 508 -407
rect 450 -447 462 -413
rect 496 -447 508 -413
rect 450 -453 508 -447
rect 941 -413 999 -407
rect 941 -447 953 -413
rect 987 -447 999 -413
rect 941 -453 999 -447
rect 462 -494 496 -453
rect 954 -494 989 -453
rect 456 -506 590 -494
rect 860 -506 994 -494
rect 443 -682 453 -506
rect 505 -682 590 -506
rect 687 -682 697 -506
rect 753 -682 763 -506
rect 860 -682 943 -506
rect 999 -682 1009 -506
rect 456 -694 590 -682
rect 860 -694 994 -682
rect 602 -784 612 -732
rect 680 -784 690 -732
rect 779 -812 831 -775
rect 619 -864 830 -812
rect 619 -898 673 -864
rect 450 -906 508 -900
rect 450 -940 462 -906
rect 496 -940 508 -906
rect 450 -946 508 -940
rect 462 -987 496 -946
rect 616 -947 676 -898
rect 760 -949 770 -897
rect 838 -949 848 -897
rect 942 -906 1000 -900
rect 942 -940 954 -906
rect 988 -940 1000 -906
rect 942 -946 1000 -940
rect 954 -987 988 -946
rect 456 -1187 590 -987
rect 860 -999 994 -987
rect 687 -1175 697 -999
rect 753 -1175 763 -999
rect 860 -1175 901 -999
rect 953 -1175 994 -999
rect 860 -1187 994 -1175
rect 495 -1435 551 -1187
rect 495 -1491 943 -1435
rect 999 -1491 1009 -1435
<< via1 >>
rect 941 748 997 804
rect 697 302 753 478
rect 901 302 953 478
rect 770 200 838 252
rect 612 36 680 88
rect 453 -190 505 -14
rect 697 -190 753 -14
rect 943 -190 999 -14
rect 453 -682 505 -506
rect 697 -682 753 -506
rect 943 -682 999 -506
rect 612 -784 680 -732
rect 770 -949 838 -897
rect 697 -1175 753 -999
rect 901 -1175 953 -999
rect 943 -1491 999 -1435
<< metal2 >>
rect 941 804 997 814
rect 941 739 997 748
rect 955 738 997 739
rect 451 632 953 684
rect 451 -4 503 632
rect 697 478 753 488
rect 697 292 753 302
rect 901 478 953 632
rect 901 292 953 302
rect 770 252 838 262
rect 770 190 838 200
rect 778 162 830 190
rect 620 129 830 162
rect 620 98 672 129
rect 612 88 680 98
rect 612 26 680 36
rect 451 -14 505 -4
rect 451 -190 453 -14
rect 451 -200 505 -190
rect 697 -14 753 -4
rect 697 -200 753 -190
rect 943 -14 999 -4
rect 943 -200 999 -190
rect 451 -496 503 -200
rect 451 -506 505 -496
rect 451 -682 453 -506
rect 451 -692 505 -682
rect 697 -506 753 -496
rect 697 -692 753 -682
rect 943 -506 999 -496
rect 943 -692 999 -682
rect 451 -1326 503 -692
rect 612 -732 680 -722
rect 612 -794 680 -784
rect 619 -822 671 -794
rect 619 -855 831 -822
rect 779 -887 831 -855
rect 770 -897 838 -887
rect 770 -959 838 -949
rect 697 -999 753 -989
rect 697 -1185 753 -1175
rect 901 -999 953 -989
rect 901 -1326 953 -1175
rect 451 -1378 953 -1326
rect 943 -1433 999 -1425
rect 941 -1435 1001 -1433
rect 941 -1491 943 -1435
rect 999 -1491 1001 -1435
rect 941 -1493 1001 -1491
rect 943 -1501 999 -1493
<< via2 >>
rect 941 748 997 804
rect 697 302 753 478
rect 697 -190 753 -14
rect 943 -190 999 -14
rect 697 -682 753 -506
rect 943 -682 999 -506
rect 697 -1175 753 -999
rect 943 -1491 999 -1435
<< metal3 >>
rect 931 804 1007 809
rect 931 748 941 804
rect 997 748 1007 804
rect 931 743 1007 748
rect 687 478 763 483
rect 687 302 697 478
rect 753 302 763 478
rect 687 297 763 302
rect 694 -9 755 297
rect 941 -9 1001 743
rect 687 -14 763 -9
rect 687 -190 697 -14
rect 753 -190 763 -14
rect 687 -195 763 -190
rect 933 -14 1009 -9
rect 933 -190 943 -14
rect 999 -190 1009 -14
rect 933 -195 1009 -190
rect 694 -501 755 -195
rect 941 -501 1001 -195
rect 687 -506 763 -501
rect 687 -682 697 -506
rect 753 -682 763 -506
rect 687 -687 763 -682
rect 933 -506 1009 -501
rect 933 -682 943 -506
rect 999 -682 1009 -506
rect 933 -687 1009 -682
rect 694 -994 755 -687
rect 687 -999 763 -994
rect 687 -1175 697 -999
rect 753 -1175 763 -999
rect 687 -1180 763 -1175
rect 694 -1186 755 -1180
rect 941 -1430 1001 -687
rect 933 -1435 1009 -1430
rect 933 -1491 943 -1435
rect 999 -1491 1009 -1435
rect 933 -1496 1009 -1491
rect 941 -1497 1001 -1496
use sky130_fd_pr__pfet_01v8_2XUZHN  sky130_fd_pr__pfet_01v8_2XUZHN_0
timestamp 1729189057
transform 1 0 927 0 1 390
box -109 -162 109 162
use sky130_fd_pr__pfet_01v8_2XUZHN  sky130_fd_pr__pfet_01v8_2XUZHN_1
timestamp 1729189057
transform 1 0 523 0 1 390
box -109 -162 109 162
use sky130_fd_pr__pfet_01v8_2XUZHN  sky130_fd_pr__pfet_01v8_2XUZHN_2
timestamp 1729189057
transform 1 0 523 0 1 -102
box -109 -162 109 162
use sky130_fd_pr__pfet_01v8_2XUZHN  sky130_fd_pr__pfet_01v8_2XUZHN_3
timestamp 1729189057
transform 1 0 927 0 1 -102
box -109 -162 109 162
use sky130_fd_pr__pfet_01v8_2XUZHN  sky130_fd_pr__pfet_01v8_2XUZHN_4
timestamp 1729189057
transform 1 0 523 0 1 -594
box -109 -162 109 162
use sky130_fd_pr__pfet_01v8_2XUZHN  sky130_fd_pr__pfet_01v8_2XUZHN_5
timestamp 1729189057
transform 1 0 927 0 1 -594
box -109 -162 109 162
use sky130_fd_pr__pfet_01v8_2XUZHN  sky130_fd_pr__pfet_01v8_2XUZHN_6
timestamp 1729189057
transform 1 0 523 0 1 -1087
box -109 -162 109 162
use sky130_fd_pr__pfet_01v8_2XUZHN  sky130_fd_pr__pfet_01v8_2XUZHN_7
timestamp 1729189057
transform 1 0 927 0 1 -1087
box -109 -162 109 162
use sky130_fd_pr__pfet_01v8_VQXXLL  sky130_fd_pr__pfet_01v8_VQXXLL_0
timestamp 1729189057
transform 1 0 725 0 1 -1087
box -223 -200 223 200
use sky130_fd_pr__pfet_01v8_VQXXLL  sky130_fd_pr__pfet_01v8_VQXXLL_1
timestamp 1729189057
transform 1 0 725 0 1 -594
box -223 -200 223 200
use sky130_fd_pr__pfet_01v8_VQXXLL  sky130_fd_pr__pfet_01v8_VQXXLL_2
timestamp 1729189057
transform 1 0 725 0 1 -102
box -223 -200 223 200
use sky130_fd_pr__pfet_01v8_VQXXLL  sky130_fd_pr__pfet_01v8_VQXXLL_3
timestamp 1729189057
transform 1 0 725 0 1 390
box -223 -200 223 200
<< labels >>
flabel viali 655 861 655 861 0 FreeSans 480 0 0 0 VDD
port 0 nsew
flabel metal1 644 184 644 184 0 FreeSans 480 0 0 0 VIP
port 3 nsew
flabel metal2 648 110 648 110 0 FreeSans 480 0 0 0 VIN
port 4 nsew
flabel metal3 724 38 724 38 0 FreeSans 480 0 0 0 D5
port 5 nsew
flabel metal2 612 652 612 652 0 FreeSans 480 0 0 0 D6
port 1 nsew
flabel metal3 974 710 974 710 0 FreeSans 480 0 0 0 OUT
port 2 nsew
<< end >>
