magic
tech sky130A
magscale 1 2
timestamp 1729182859
<< error_p >>
rect -269 181 -205 187
rect -111 181 -47 187
rect 47 181 111 187
rect 205 181 269 187
rect -269 147 -257 181
rect -111 147 -99 181
rect 47 147 59 181
rect 205 147 217 181
rect -269 141 -205 147
rect -111 141 -47 147
rect 47 141 111 147
rect 205 141 269 147
rect -269 -147 -205 -141
rect -111 -147 -47 -141
rect 47 -147 111 -141
rect 205 -147 269 -141
rect -269 -181 -257 -147
rect -111 -181 -99 -147
rect 47 -181 59 -147
rect 205 -181 217 -147
rect -269 -187 -205 -181
rect -111 -187 -47 -181
rect 47 -187 111 -181
rect 205 -187 269 -181
<< nwell >>
rect -381 -200 381 200
<< pmos >>
rect -287 -100 -187 100
rect -129 -100 -29 100
rect 29 -100 129 100
rect 187 -100 287 100
<< pdiff >>
rect -345 88 -287 100
rect -345 -88 -333 88
rect -299 -88 -287 88
rect -345 -100 -287 -88
rect -187 88 -129 100
rect -187 -88 -175 88
rect -141 -88 -129 88
rect -187 -100 -129 -88
rect -29 88 29 100
rect -29 -88 -17 88
rect 17 -88 29 88
rect -29 -100 29 -88
rect 129 88 187 100
rect 129 -88 141 88
rect 175 -88 187 88
rect 129 -100 187 -88
rect 287 88 345 100
rect 287 -88 299 88
rect 333 -88 345 88
rect 287 -100 345 -88
<< pdiffc >>
rect -333 -88 -299 88
rect -175 -88 -141 88
rect -17 -88 17 88
rect 141 -88 175 88
rect 299 -88 333 88
<< poly >>
rect -287 181 -187 197
rect -287 147 -271 181
rect -203 147 -187 181
rect -287 100 -187 147
rect -129 181 -29 197
rect -129 147 -113 181
rect -45 147 -29 181
rect -129 100 -29 147
rect 29 181 129 197
rect 29 147 45 181
rect 113 147 129 181
rect 29 100 129 147
rect 187 181 287 197
rect 187 147 203 181
rect 271 147 287 181
rect 187 100 287 147
rect -287 -147 -187 -100
rect -287 -181 -271 -147
rect -203 -181 -187 -147
rect -287 -197 -187 -181
rect -129 -147 -29 -100
rect -129 -181 -113 -147
rect -45 -181 -29 -147
rect -129 -197 -29 -181
rect 29 -147 129 -100
rect 29 -181 45 -147
rect 113 -181 129 -147
rect 29 -197 129 -181
rect 187 -147 287 -100
rect 187 -181 203 -147
rect 271 -181 287 -147
rect 187 -197 287 -181
<< polycont >>
rect -271 147 -203 181
rect -113 147 -45 181
rect 45 147 113 181
rect 203 147 271 181
rect -271 -181 -203 -147
rect -113 -181 -45 -147
rect 45 -181 113 -147
rect 203 -181 271 -147
<< locali >>
rect -287 147 -271 181
rect -203 147 -187 181
rect -129 147 -113 181
rect -45 147 -29 181
rect 29 147 45 181
rect 113 147 129 181
rect 187 147 203 181
rect 271 147 287 181
rect -333 88 -299 104
rect -333 -104 -299 -88
rect -175 88 -141 104
rect -175 -104 -141 -88
rect -17 88 17 104
rect -17 -104 17 -88
rect 141 88 175 104
rect 141 -104 175 -88
rect 299 88 333 104
rect 299 -104 333 -88
rect -287 -181 -271 -147
rect -203 -181 -187 -147
rect -129 -181 -113 -147
rect -45 -181 -29 -147
rect 29 -181 45 -147
rect 113 -181 129 -147
rect 187 -181 203 -147
rect 271 -181 287 -147
<< viali >>
rect -257 147 -217 181
rect -99 147 -59 181
rect 59 147 99 181
rect 217 147 257 181
rect -333 -88 -299 88
rect -175 -88 -141 88
rect -17 -88 17 88
rect 141 -88 175 88
rect 299 -88 333 88
rect -257 -181 -217 -147
rect -99 -181 -59 -147
rect 59 -181 99 -147
rect 217 -181 257 -147
<< metal1 >>
rect -269 181 -205 187
rect -269 147 -257 181
rect -217 147 -205 181
rect -269 141 -205 147
rect -111 181 -47 187
rect -111 147 -99 181
rect -59 147 -47 181
rect -111 141 -47 147
rect 47 181 111 187
rect 47 147 59 181
rect 99 147 111 181
rect 47 141 111 147
rect 205 181 269 187
rect 205 147 217 181
rect 257 147 269 181
rect 205 141 269 147
rect -339 88 -293 100
rect -339 -88 -333 88
rect -299 -88 -293 88
rect -339 -100 -293 -88
rect -181 88 -135 100
rect -181 -88 -175 88
rect -141 -88 -135 88
rect -181 -100 -135 -88
rect -23 88 23 100
rect -23 -88 -17 88
rect 17 -88 23 88
rect -23 -100 23 -88
rect 135 88 181 100
rect 135 -88 141 88
rect 175 -88 181 88
rect 135 -100 181 -88
rect 293 88 339 100
rect 293 -88 299 88
rect 333 -88 339 88
rect 293 -100 339 -88
rect -269 -147 -205 -141
rect -269 -181 -257 -147
rect -217 -181 -205 -147
rect -269 -187 -205 -181
rect -111 -147 -47 -141
rect -111 -181 -99 -147
rect -59 -181 -47 -147
rect -111 -187 -47 -181
rect 47 -147 111 -141
rect 47 -181 59 -147
rect 99 -181 111 -147
rect 47 -187 111 -181
rect 205 -147 269 -141
rect 205 -181 217 -147
rect 257 -181 269 -147
rect 205 -187 269 -181
<< properties >>
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 1 l 0.5 m 1 nf 4 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 60 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
