* PEX produced on Fri Oct 18 15:01:37 WIB 2024 using ./iic-pex.sh with m=3 and s=1
* NGSPICE file created from opamp.ext - technology: sky130A

.subckt opamp OUT GND VIN VIP RS VDD
X0 VDD.t22 VDD.t20 VDD.t21 VDD.t1 sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0 ps=0 w=2 l=0.15
X1 VDD.t19 VDD.t18 VDD.t19 VDD.t4 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.29 as=0 ps=0 w=2 l=0.15
X2 VDD.t13 pmoscs_0.D2.t17 pmosdif_0.D5.t2 VDD.t8 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X3 VDD.t9 pmoscs_0.D2.t13 pmoscs_0.D2.t14 VDD.t8 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X4 GND.t13 pmoscs_0.D1.t2 pmoscs_0.D1.t3 GND.t12 sky130_fd_pr__nfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=1
X5 pmoscs_0.D1.t14 pmoscs_0.D1.t12 pmoscs_0.D1.t13 GND.t0 sky130_fd_pr__nfet_01v8 ad=0.58 pd=4.58 as=0 ps=0 w=2 l=0.15
X6 OUT.t22 pmosdif_0.D6.t27 GND.t16 GND.t14 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.8
X7 pmosdif_0.D5.t0 VIP.t0 OUT.t0 VDD.t0 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X8 pmoscs_0.D1.t11 pmoscs_0.D1.t9 pmoscs_0.D1.t10 GND.t1 sky130_fd_pr__nfet_01v8 ad=0.58 pd=4.58 as=0 ps=0 w=2 l=0.15
X9 OUT.t16 OUT.t14 OUT.t15 GND.t7 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.15
X10 pmosdif_0.D6.t26 pmosdif_0.D6.t25 pmosdif_0.D6.t26 GND.t2 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0 ps=0 w=1 l=0.15
X11 pmoscs_0.D2.t10 pmoscs_0.D2.t9 pmoscs_0.D2.t10 VDD.t4 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.29 as=0 ps=0 w=2 l=0.15
X12 GND.t19 pmosdif_0.D6.t28 OUT.t21 GND.t5 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.8
X13 OUT.t13 OUT.t12 OUT.t13 VDD.t2 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0 ps=0 w=1 l=0.15
X14 VDD.t11 pmoscs_0.D2.t18 pmoscs_0.D1.t1 VDD.t8 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X15 OUT.t20 pmosdif_0.D6.t29 GND.t18 GND.t8 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.8
X16 VDD.t17 VDD.t16 VDD.t17 VDD.t8 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.29 as=0 ps=0 w=2 l=1
X17 RS.t1 pmoscs_0.D1.t17 pmoscs_0.D2.t15 GND.t12 sky130_fd_pr__nfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=1
X18 pmoscs_0.D1.t8 pmoscs_0.D1.t7 pmoscs_0.D1.t8 VDD.t4 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.29 as=0 ps=0 w=2 l=0.15
X19 pmoscs_0.D2.t8 pmoscs_0.D2.t6 pmoscs_0.D2.t7 GND.t1 sky130_fd_pr__nfet_01v8 ad=0.58 pd=4.58 as=0 ps=0 w=2 l=0.15
X20 OUT.t11 OUT.t9 OUT.t10 VDD.t3 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.15
X21 pmosdif_0.D6.t24 pmosdif_0.D6.t22 pmosdif_0.D6.t23 VDD.t3 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.15
X22 pmosdif_0.D6.t2 VIN.t0 pmosdif_0.D5.t7 VDD.t5 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X23 pmosdif_0.D5.t3 VIN.t1 pmosdif_0.D6.t0 VDD.t0 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X24 OUT.t8 OUT.t7 OUT.t8 GND.t2 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0 ps=0 w=1 l=0.15
X25 GND.t4 pmosdif_0.D6.t10 pmosdif_0.D6.t11 GND.t3 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.8
X26 pmosdif_0.D5.t14 pmosdif_0.D5.t13 pmosdif_0.D5.t14 VDD.t4 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.29 as=0 ps=0 w=2 l=0.15
X27 GND.t6 pmosdif_0.D6.t8 pmosdif_0.D6.t9 GND.t5 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.8
X28 pmoscs_0.D2.t16 pmoscs_0.D1.t18 RS.t0 GND.t10 sky130_fd_pr__nfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=1
X29 pmosdif_0.D6.t7 pmosdif_0.D6.t6 GND.t9 GND.t8 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.8
X30 OUT.t6 OUT.t5 OUT.t6 VDD.t2 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0 ps=0 w=1 l=0.15
X31 OUT.t4 OUT.t2 OUT.t3 VDD.t3 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.15
X32 pmosdif_0.D6.t21 pmosdif_0.D6.t19 pmosdif_0.D6.t20 VDD.t3 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.15
X33 OUT.t1 VIP.t1 pmosdif_0.D5.t4 VDD.t5 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X34 pmosdif_0.D5.t5 VIN.t2 pmosdif_0.D6.t1 VDD.t0 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X35 pmoscs_0.D1.t16 pmoscs_0.D1.t15 GND.t11 GND.t10 sky130_fd_pr__nfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=1
X36 OUT.t17 VIP.t2 pmosdif_0.D5.t6 VDD.t5 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X37 GND.t17 pmosdif_0.D6.t30 OUT.t19 GND.t3 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.8
X38 pmosdif_0.D6.t18 pmosdif_0.D6.t17 pmosdif_0.D6.t18 VDD.t2 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0 ps=0 w=1 l=0.15
X39 pmoscs_0.D1.t0 pmoscs_0.D2.t19 VDD.t12 VDD.t6 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X40 VDD.t15 VDD.t14 VDD.t15 VDD.t6 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.29 as=0 ps=0 w=2 l=1
X41 pmosdif_0.D6.t16 pmosdif_0.D6.t14 pmosdif_0.D6.t15 GND.t7 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.15
X42 pmosdif_0.D6.t5 pmosdif_0.D6.t4 GND.t15 GND.t14 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.8
X43 pmosdif_0.D5.t12 pmosdif_0.D5.t10 pmosdif_0.D5.t11 VDD.t1 sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0 ps=0 w=2 l=0.15
X44 pmoscs_0.D2.t5 pmoscs_0.D2.t3 pmoscs_0.D2.t4 VDD.t1 sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0 ps=0 w=2 l=0.15
X45 pmosdif_0.D5.t9 VIP.t3 OUT.t18 VDD.t0 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X46 pmosdif_0.D6.t13 pmosdif_0.D6.t12 pmosdif_0.D6.t13 VDD.t2 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0 ps=0 w=1 l=0.15
X47 pmoscs_0.D2.t2 pmoscs_0.D2.t0 pmoscs_0.D2.t1 GND.t0 sky130_fd_pr__nfet_01v8 ad=0.58 pd=4.58 as=0 ps=0 w=2 l=0.15
X48 pmosdif_0.D6.t3 VIN.t3 pmosdif_0.D5.t8 VDD.t5 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X49 pmoscs_0.D1.t6 pmoscs_0.D1.t4 pmoscs_0.D1.t5 VDD.t1 sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0 ps=0 w=2 l=0.15
X50 pmoscs_0.D2.t12 pmoscs_0.D2.t11 VDD.t7 VDD.t6 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X51 pmosdif_0.D5.t1 pmoscs_0.D2.t20 VDD.t10 VDD.t6 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
R0 VDD.n8 VDD.n7 39566.1
R1 VDD.n40 VDD.n39 23430.6
R2 VDD.n42 VDD.n15 6391.76
R3 VDD.n38 VDD.n15 6388.23
R4 VDD.n42 VDD.n14 6384.71
R5 VDD.n38 VDD.n14 6381.18
R6 VDD.n5 VDD.n2 5403.53
R7 VDD.n9 VDD.n2 5403.53
R8 VDD.n5 VDD.n3 5403.53
R9 VDD.n9 VDD.n3 5403.53
R10 VDD.n43 VDD.n13 681.788
R11 VDD.n37 VDD.n12 680.659
R12 VDD.n10 VDD.n1 576.378
R13 VDD.n4 VDD.n1 576.378
R14 VDD.n4 VDD.n0 575.914
R15 VDD.n34 VDD.t20 555.769
R16 VDD.n20 VDD.t18 555.274
R17 VDD.n11 VDD.n10 551.907
R18 VDD.n44 VDD.n12 551.337
R19 VDD.n36 VDD.n13 550.777
R20 VDD.n23 VDD.t14 144.274
R21 VDD.n16 VDD.t16 144.274
R22 VDD.n37 VDD.n36 130.636
R23 VDD.n44 VDD.n43 129.323
R24 VDD.n21 VDD.t19 111.784
R25 VDD.n33 VDD.t22 111.784
R26 VDD.n30 VDD.n29 100.016
R27 VDD.n24 VDD.n17 100.013
R28 VDD.n22 VDD.n19 99.3605
R29 VDD.n26 VDD.n25 99.3605
R30 VDD.n28 VDD.n27 99.3605
R31 VDD.n32 VDD.n31 99.3605
R32 VDD.n21 VDD.n20 96.2857
R33 VDD.n34 VDD.n33 96.2857
R34 VDD.t2 VDD.n5 59.9871
R35 VDD.t6 VDD.t4 57.3252
R36 VDD.t8 VDD.t1 57.3252
R37 VDD.n8 VDD.t3 55.3035
R38 VDD.t4 VDD.n14 52.4595
R39 VDD.t1 VDD.n39 47.7159
R40 VDD.t5 VDD.t2 46.5914
R41 VDD.t0 VDD.t3 46.5914
R42 VDD.n41 VDD.t6 42.4142
R43 VDD.n40 VDD.t8 42.4142
R44 VDD.n6 VDD.t5 30.3035
R45 VDD.n7 VDD.t0 29.1672
R46 VDD.n11 VDD.n0 22.6748
R47 VDD.n3 VDD.n1 20.5561
R48 VDD.n6 VDD.n3 20.5561
R49 VDD.n2 VDD.n0 20.5561
R50 VDD.n6 VDD.n2 20.5561
R51 VDD.n43 VDD.n42 15.4172
R52 VDD.n42 VDD.n41 15.4172
R53 VDD.n38 VDD.n37 15.4172
R54 VDD.n41 VDD.n38 15.4172
R55 VDD.t19 VDD.n19 14.283
R56 VDD.n19 VDD.t15 14.283
R57 VDD.n25 VDD.t7 14.283
R58 VDD.n25 VDD.t11 14.283
R59 VDD.n27 VDD.t12 14.283
R60 VDD.n27 VDD.t9 14.283
R61 VDD.n30 VDD.t10 14.283
R62 VDD.t17 VDD.n30 14.283
R63 VDD.n31 VDD.t17 14.283
R64 VDD.n31 VDD.t21 14.283
R65 VDD.t15 VDD.n17 14.283
R66 VDD.n17 VDD.t13 14.283
R67 VDD.n36 VDD.n35 9.47742
R68 VDD.n35 VDD.n34 9.3005
R69 VDD.n20 VDD.n18 9.3005
R70 VDD.n45 VDD.n44 9.3005
R71 VDD.n10 VDD.n9 5.44168
R72 VDD.n9 VDD.n8 5.44168
R73 VDD.n5 VDD.n4 5.44168
R74 VDD.n14 VDD.n12 4.74409
R75 VDD.n15 VDD.n13 4.74409
R76 VDD.n39 VDD.n15 4.74409
R77 VDD.n46 VDD.n45 3.91791
R78 VDD VDD.n11 3.11912
R79 VDD.n46 VDD 2.02187
R80 VDD.n28 VDD.n26 1.88909
R81 VDD.n33 VDD.n32 1.8605
R82 VDD.n22 VDD.n21 1.8605
R83 VDD VDD.n47 1.48407
R84 VDD.n29 VDD.n28 1.1092
R85 VDD.n26 VDD.n24 1.10648
R86 VDD.n41 VDD.n40 0.663214
R87 VDD.n32 VDD.n16 0.649024
R88 VDD.n23 VDD.n22 0.629776
R89 VDD.n22 VDD.n18 0.387371
R90 VDD.n7 VDD.n6 0.379288
R91 VDD.n29 VDD.n16 0.351043
R92 VDD.n35 VDD.n32 0.348049
R93 VDD.n24 VDD.n23 0.336438
R94 VDD VDD.n46 0.164562
R95 VDD.n18 VDD 0.119922
R96 VDD.n45 VDD 0.0849275
R97 pmoscs_0.D2.n6 pmoscs_0.D2.t3 563.553
R98 pmoscs_0.D2.n4 pmoscs_0.D2.t9 556.88
R99 pmoscs_0.D2.n2 pmoscs_0.D2.t0 549.227
R100 pmoscs_0.D2.n17 pmoscs_0.D2.t6 540.813
R101 pmoscs_0.D2.t18 pmoscs_0.D2.t17 167.495
R102 pmoscs_0.D2.t19 pmoscs_0.D2.t20 167.495
R103 pmoscs_0.D2.n16 pmoscs_0.D2.t11 144.931
R104 pmoscs_0.D2.n6 pmoscs_0.D2.t5 113.382
R105 pmoscs_0.D2.t10 pmoscs_0.D2.n5 111.784
R106 pmoscs_0.D2.n8 pmoscs_0.D2.n7 99.3605
R107 pmoscs_0.D2.n15 pmoscs_0.D2.n14 99.3605
R108 pmoscs_0.D2.n17 pmoscs_0.D2.n3 92.8975
R109 pmoscs_0.D2.n10 pmoscs_0.D2.n9 85.4606
R110 pmoscs_0.D2 pmoscs_0.D2.n13 85.4606
R111 pmoscs_0.D2.n11 pmoscs_0.D2.t18 83.8685
R112 pmoscs_0.D2.n12 pmoscs_0.D2.t19 83.6275
R113 pmoscs_0.D2.n5 pmoscs_0.D2.n4 70.4685
R114 pmoscs_0.D2.n10 pmoscs_0.D2.t13 63.6245
R115 pmoscs_0.D2.n13 pmoscs_0.D2.t11 63.6245
R116 pmoscs_0.D2.n1 pmoscs_0.D2.t16 41.4116
R117 pmoscs_0.D2.n0 pmoscs_0.D2.t15 41.4116
R118 pmoscs_0.D2.n1 pmoscs_0.D2.t2 41.3938
R119 pmoscs_0.D2.n0 pmoscs_0.D2.t7 41.3938
R120 pmoscs_0.D2.n2 pmoscs_0.D2.t1 41.1927
R121 pmoscs_0.D2.n3 pmoscs_0.D2.t8 39.5338
R122 pmoscs_0.D2.n12 pmoscs_0.D2.n11 27.6797
R123 pmoscs_0.D2.n13 pmoscs_0.D2.n12 20.2445
R124 pmoscs_0.D2.n11 pmoscs_0.D2.n10 20.0035
R125 pmoscs_0.D2.n7 pmoscs_0.D2.t14 14.283
R126 pmoscs_0.D2.n7 pmoscs_0.D2.t4 14.283
R127 pmoscs_0.D2.n14 pmoscs_0.D2.t10 14.283
R128 pmoscs_0.D2.n14 pmoscs_0.D2.t12 14.283
R129 pmoscs_0.D2.n18 pmoscs_0.D2.n17 9.3005
R130 pmoscs_0.D2.n16 pmoscs_0.D2.n4 9.3005
R131 pmoscs_0.D2.n16 pmoscs_0.D2.n15 5.8147
R132 pmoscs_0.D2 pmoscs_0.D2.n0 2.24018
R133 pmoscs_0.D2.n0 pmoscs_0.D2.n3 1.8605
R134 pmoscs_0.D2.n15 pmoscs_0.D2.n5 1.8605
R135 pmoscs_0.D2 pmoscs_0.D2.n1 1.5981
R136 pmoscs_0.D2 pmoscs_0.D2.n9 1.50561
R137 pmoscs_0.D2.n9 pmoscs_0.D2.n8 1.38512
R138 pmoscs_0.D2.n15 pmoscs_0.D2 1.3734
R139 pmoscs_0.D2.n18 pmoscs_0.D2.n16 1.0364
R140 pmoscs_0.D2.n8 pmoscs_0.D2.n6 0.21948
R141 pmoscs_0.D2.n1 pmoscs_0.D2.n2 0.214768
R142 pmoscs_0.D2.n0 pmoscs_0.D2.n18 0.132769
R143 pmosdif_0.D5.n2 pmosdif_0.D5.t10 564.03
R144 pmosdif_0.D5.n7 pmosdif_0.D5.t13 549.005
R145 pmosdif_0.D5.n6 pmosdif_0.D5.n4 203.958
R146 pmosdif_0.D5 pmosdif_0.D5.n3 203.863
R147 pmosdif_0.D5.n6 pmosdif_0.D5.n5 203.606
R148 pmosdif_0.D5 pmosdif_0.D5.n13 203.606
R149 pmosdif_0.D5.t14 pmosdif_0.D5.n7 113.374
R150 pmosdif_0.D5.n1 pmosdif_0.D5.n10 99.3605
R151 pmosdif_0.D5.n9 pmosdif_0.D5.n8 99.3605
R152 pmosdif_0.D5.t12 pmosdif_0.D5.n2 113.343
R153 pmosdif_0.D5.n5 pmosdif_0.D5.t6 28.5655
R154 pmosdif_0.D5.n5 pmosdif_0.D5.t5 28.5655
R155 pmosdif_0.D5.n4 pmosdif_0.D5.t8 28.5655
R156 pmosdif_0.D5.n4 pmosdif_0.D5.t9 28.5655
R157 pmosdif_0.D5.n13 pmosdif_0.D5.t4 28.5655
R158 pmosdif_0.D5.n13 pmosdif_0.D5.t3 28.5655
R159 pmosdif_0.D5.n3 pmosdif_0.D5.t7 28.5655
R160 pmosdif_0.D5.n3 pmosdif_0.D5.t0 28.5655
R161 pmosdif_0.D5.n10 pmosdif_0.D5.t2 14.283
R162 pmosdif_0.D5.n10 pmosdif_0.D5.t11 14.283
R163 pmosdif_0.D5.n8 pmosdif_0.D5.t14 14.283
R164 pmosdif_0.D5.n8 pmosdif_0.D5.t1 14.283
R165 pmosdif_0.D5.n12 pmosdif_0.D5.n11 10.6783
R166 pmosdif_0.D5.n11 pmosdif_0.D5 9.13431
R167 pmosdif_0.D5.n0 pmosdif_0.D5 5.6496
R168 pmosdif_0.D5.n1 pmosdif_0.D5.n2 0.25683
R169 pmosdif_0.D5.n11 pmosdif_0.D5.n1 1.58133
R170 pmosdif_0.D5.n12 pmosdif_0.D5.n9 1.57893
R171 pmosdif_0.D5 pmosdif_0.D5.n12 1.39782
R172 pmosdif_0.D5.n9 pmosdif_0.D5.n7 0.227707
R173 pmosdif_0.D5.n0 pmosdif_0.D5.n6 0.200554
R174 pmosdif_0.D5 pmosdif_0.D5.n0 0.197969
R175 pmoscs_0.D1.n3 pmoscs_0.D1.t7 564.254
R176 pmoscs_0.D1.n6 pmoscs_0.D1.t4 563.923
R177 pmoscs_0.D1.n11 pmoscs_0.D1.t12 549.227
R178 pmoscs_0.D1.n9 pmoscs_0.D1.t9 540.813
R179 pmoscs_0.D1.t8 pmoscs_0.D1.n3 113.439
R180 pmoscs_0.D1.n6 pmoscs_0.D1.t6 113.371
R181 pmoscs_0.D1.n8 pmoscs_0.D1.n7 99.3605
R182 pmoscs_0.D1.n5 pmoscs_0.D1.n4 99.3605
R183 pmoscs_0.D1.n10 pmoscs_0.D1.n9 92.8975
R184 pmoscs_0.D1.n12 pmoscs_0.D1.n2 85.738
R185 pmoscs_0.D1 pmoscs_0.D1.n15 85.651
R186 pmoscs_0.D1.n14 pmoscs_0.D1.n13 85.4685
R187 pmoscs_0.D1.n13 pmoscs_0.D1.t18 81.2175
R188 pmoscs_0.D1.n14 pmoscs_0.D1.t17 80.9765
R189 pmoscs_0.D1.n15 pmoscs_0.D1.t2 61.4555
R190 pmoscs_0.D1.n12 pmoscs_0.D1.t15 61.4555
R191 pmoscs_0.D1.n2 pmoscs_0.D1.t16 41.3938
R192 pmoscs_0.D1.n1 pmoscs_0.D1.t10 41.3938
R193 pmoscs_0.D1.n1 pmoscs_0.D1.t3 41.3938
R194 pmoscs_0.D1.n2 pmoscs_0.D1.t14 41.3938
R195 pmoscs_0.D1.n11 pmoscs_0.D1.t13 41.1927
R196 pmoscs_0.D1.n10 pmoscs_0.D1.t11 39.5338
R197 pmoscs_0.D1.n15 pmoscs_0.D1.n14 19.7625
R198 pmoscs_0.D1.n13 pmoscs_0.D1.n12 19.5215
R199 pmoscs_0.D1.n7 pmoscs_0.D1.t1 14.283
R200 pmoscs_0.D1.n7 pmoscs_0.D1.t5 14.283
R201 pmoscs_0.D1.n4 pmoscs_0.D1.t8 14.283
R202 pmoscs_0.D1.n4 pmoscs_0.D1.t0 14.283
R203 pmoscs_0.D1.n9 pmoscs_0.D1.n0 9.3005
R204 pmoscs_0.D1.n0 pmoscs_0.D1 8.95986
R205 pmoscs_0.D1 pmoscs_0.D1.n8 2.03536
R206 pmoscs_0.D1.n1 pmoscs_0.D1.n10 1.8605
R207 pmoscs_0.D1 pmoscs_0.D1.n5 1.6418
R208 pmoscs_0.D1.n2 pmoscs_0.D1.n11 0.23258
R209 pmoscs_0.D1.n8 pmoscs_0.D1.n6 0.230482
R210 pmoscs_0.D1.n5 pmoscs_0.D1.n3 0.174465
R211 pmoscs_0.D1.n1 pmoscs_0.D1.n0 0.134277
R212 pmoscs_0.D1 pmoscs_0.D1.n1 0.0874565
R213 GND.n34 GND.n6 7903.18
R214 GND.n34 GND.n7 7903.18
R215 GND.n19 GND.n6 7880
R216 GND.n19 GND.n7 7880
R217 GND.n9 GND.n8 7486
R218 GND.n32 GND.n8 7486
R219 GND.n32 GND.n27 7486
R220 GND.n27 GND.n9 7486
R221 GND.t12 GND.n24 1471.8
R222 GND.n24 GND.n23 1348.51
R223 GND.n18 GND.n4 512
R224 GND.n28 GND.n1 486.401
R225 GND.n31 GND.n2 486.401
R226 GND.n36 GND.n35 467.627
R227 GND.n31 GND.n30 463.06
R228 GND.n18 GND.n17 388.228
R229 GND.n35 GND.n5 386.733
R230 GND.n26 GND.t12 340.382
R231 GND.n22 GND.t8 301.175
R232 GND.t2 GND.n19 296.75
R233 GND.n39 GND.n38 285.784
R234 GND.t0 GND.n20 274.443
R235 GND.t14 GND.t2 272.661
R236 GND.n33 GND.t7 249.494
R237 GND.t10 GND.n21 222.895
R238 GND.n25 GND.t1 215.659
R239 GND.t12 GND.n25 199.738
R240 GND.n21 GND.t0 192.501
R241 GND.n39 GND.n1 180.373
R242 GND.n10 GND.n5 126.204
R243 GND.n17 GND.n10 123.204
R244 GND.n11 GND.t6 83.7528
R245 GND.n11 GND.t16 83.7528
R246 GND.n12 GND.t19 83.7528
R247 GND.n12 GND.t15 83.7528
R248 GND.n13 GND.t17 83.7528
R249 GND.n13 GND.t9 83.7528
R250 GND.n14 GND.t4 83.7528
R251 GND.n14 GND.t18 83.7528
R252 GND.n20 GND.t14 80.1949
R253 GND.n36 GND.n4 44.4749
R254 GND.n34 GND.n33 43.6914
R255 GND.n3 GND.t11 41.3938
R256 GND.n29 GND.t13 41.3938
R257 GND.n35 GND.n34 36.563
R258 GND.n19 GND.n18 36.563
R259 GND.n28 GND.n8 34.4123
R260 GND.n24 GND.n8 34.4123
R261 GND.n27 GND.n2 34.4123
R262 GND.n27 GND.n26 34.4123
R263 GND.n9 GND.n1 30.79
R264 GND.n20 GND.n9 30.79
R265 GND.n32 GND.n31 30.79
R266 GND.n33 GND.n32 30.79
R267 GND.n10 GND.n7 26.5914
R268 GND.n22 GND.n7 26.5914
R269 GND.n6 GND.n4 26.5914
R270 GND.n22 GND.n6 26.5914
R271 GND.n25 GND.t3 23.9826
R272 GND.n21 GND.t5 23.8893
R273 GND.n30 GND.n28 23.3417
R274 GND.n38 GND.n2 19.577
R275 GND.n17 GND.n16 13.9688
R276 GND.n15 GND.n5 13.9664
R277 GND.n37 GND.n36 9.85556
R278 GND GND.n39 9.5966
R279 GND.n30 GND 9.49918
R280 GND.n38 GND.n37 9.3005
R281 GND.n23 GND.t10 8.68471
R282 GND.t1 GND.t7 7.12889
R283 GND.n23 GND.n22 5.34679
R284 GND.n26 GND.t8 5.34679
R285 GND.n15 GND.n14 2.78982
R286 GND GND.n12 2.65915
R287 GND.n29 GND.n3 2.01409
R288 GND.n16 GND.n15 1.59906
R289 GND GND.n0 1.29219
R290 GND.n37 GND.n3 0.957135
R291 GND GND.n29 0.726043
R292 GND.n12 GND.n11 0.708833
R293 GND.n14 GND.n13 0.708833
R294 GND.n16 GND 0.132712
R295 pmosdif_0.D6.n8 pmosdif_0.D6.t19 403.365
R296 pmosdif_0.D6.n12 pmosdif_0.D6.t22 402.632
R297 pmosdif_0.D6.n16 pmosdif_0.D6.t17 402.327
R298 pmosdif_0.D6.n6 pmosdif_0.D6.t12 402.327
R299 pmosdif_0.D6.n4 pmosdif_0.D6.t25 387.755
R300 pmosdif_0.D6.n2 pmosdif_0.D6.t14 387.755
R301 pmosdif_0.D6.t18 pmosdif_0.D6.n16 227.308
R302 pmosdif_0.D6.n6 pmosdif_0.D6.t13 227.308
R303 pmosdif_0.D6.n12 pmosdif_0.D6.t24 227.285
R304 pmosdif_0.D6.n8 pmosdif_0.D6.t21 227.282
R305 pmosdif_0.D6.n18 pmosdif_0.D6.n17 199.65
R306 pmosdif_0.D6.n14 pmosdif_0.D6.n13 199.65
R307 pmosdif_0.D6.n10 pmosdif_0.D6.n9 199.65
R308 pmosdif_0.D6.n7 pmosdif_0.D6.n5 199.65
R309 pmosdif_0.D6 pmosdif_0.D6.t10 129.675
R310 pmosdif_0.D6.n24 pmosdif_0.D6.t4 129.675
R311 pmosdif_0.D6 pmosdif_0.D6.t30 129.673
R312 pmosdif_0.D6.n24 pmosdif_0.D6.t27 129.673
R313 pmosdif_0.D6.n1 pmosdif_0.D6.t29 129.595
R314 pmosdif_0.D6.n23 pmosdif_0.D6.t28 129.595
R315 pmosdif_0.D6.n21 pmosdif_0.D6.t8 127.766
R316 pmosdif_0.D6.n21 pmosdif_0.D6.t6 127.766
R317 pmosdif_0.D6.n20 pmosdif_0.D6.t7 83.7172
R318 pmosdif_0.D6.n20 pmosdif_0.D6.t9 83.7172
R319 pmosdif_0.D6.t26 pmosdif_0.D6.n4 82.7662
R320 pmosdif_0.D6.n2 pmosdif_0.D6.t16 82.7662
R321 pmosdif_0.D6.n0 pmosdif_0.D6.n3 66.3172
R322 pmosdif_0.D6.n27 pmosdif_0.D6.n26 66.3172
R323 pmosdif_0.D6.n17 pmosdif_0.D6.t18 28.5655
R324 pmosdif_0.D6.n17 pmosdif_0.D6.t3 28.5655
R325 pmosdif_0.D6.n13 pmosdif_0.D6.t1 28.5655
R326 pmosdif_0.D6.n13 pmosdif_0.D6.t23 28.5655
R327 pmosdif_0.D6.n9 pmosdif_0.D6.t0 28.5655
R328 pmosdif_0.D6.n9 pmosdif_0.D6.t20 28.5655
R329 pmosdif_0.D6.t13 pmosdif_0.D6.n5 28.5655
R330 pmosdif_0.D6.n5 pmosdif_0.D6.t2 28.5655
R331 pmosdif_0.D6.n3 pmosdif_0.D6.t11 17.4005
R332 pmosdif_0.D6.n3 pmosdif_0.D6.t15 17.4005
R333 pmosdif_0.D6.n26 pmosdif_0.D6.t26 17.4005
R334 pmosdif_0.D6.n26 pmosdif_0.D6.t5 17.4005
R335 pmosdif_0.D6.n19 pmosdif_0.D6.n18 4.6904
R336 pmosdif_0.D6.n22 pmosdif_0.D6.n21 4.6279
R337 pmosdif_0.D6.n0 pmosdif_0.D6.n27 3.91489
R338 pmosdif_0.D6 pmosdif_0.D6.n7 3.58944
R339 pmosdif_0.D6 pmosdif_0.D6.n0 2.97406
R340 pmosdif_0.D6.n27 pmosdif_0.D6.n25 2.75531
R341 pmosdif_0.D6.n11 pmosdif_0.D6.n10 2.2505
R342 pmosdif_0.D6.n15 pmosdif_0.D6.n14 2.2505
R343 pmosdif_0.D6.n11 pmosdif_0.D6 2.08072
R344 pmosdif_0.D6.n15 pmosdif_0.D6.n11 1.16574
R345 pmosdif_0.D6.n25 pmosdif_0.D6.n19 0.925981
R346 pmosdif_0.D6.n19 pmosdif_0.D6.n15 0.842737
R347 pmosdif_0.D6.n0 pmosdif_0.D6.n2 0.643096
R348 pmosdif_0.D6.n27 pmosdif_0.D6.n4 0.64123
R349 pmosdif_0.D6.n10 pmosdif_0.D6.n8 0.639383
R350 pmosdif_0.D6.n14 pmosdif_0.D6.n12 0.637315
R351 pmosdif_0.D6.n18 pmosdif_0.D6.n16 0.61309
R352 pmosdif_0.D6.n7 pmosdif_0.D6.n6 0.61309
R353 pmosdif_0.D6.n24 pmosdif_0.D6.n23 0.546829
R354 pmosdif_0.D6 pmosdif_0.D6.n1 0.546829
R355 pmosdif_0.D6.n23 pmosdif_0.D6.n22 0.301636
R356 pmosdif_0.D6.n22 pmosdif_0.D6.n1 0.301636
R357 pmosdif_0.D6.n25 pmosdif_0.D6.n24 0.214442
R358 pmosdif_0.D6.n21 pmosdif_0.D6.n20 0.155708
R359 OUT.n3 OUT.t12 404.25
R360 OUT.n11 OUT.t2 402.327
R361 OUT.n7 OUT.t5 401.959
R362 OUT.n1 OUT.t9 401.649
R363 OUT.n16 OUT.t7 387.752
R364 OUT.n19 OUT.t14 372.909
R365 OUT.n1 OUT.t11 227.335
R366 OUT.t6 OUT.n7 227.314
R367 OUT.n11 OUT.t4 227.308
R368 OUT.t13 OUT.n3 227.29
R369 OUT.n13 OUT.n12 199.65
R370 OUT.n9 OUT.n8 199.65
R371 OUT.n5 OUT.n4 199.65
R372 OUT.n2 OUT.n0 199.65
R373 OUT.n22 OUT.t20 83.7528
R374 OUT.n22 OUT.t21 83.7528
R375 OUT.n19 OUT.t16 82.7664
R376 OUT.n16 OUT.t8 82.7664
R377 OUT.n20 OUT.n18 66.3172
R378 OUT.n17 OUT.n15 66.3172
R379 OUT.n12 OUT.t18 28.5655
R380 OUT.n12 OUT.t3 28.5655
R381 OUT.n8 OUT.t6 28.5655
R382 OUT.n8 OUT.t17 28.5655
R383 OUT.n4 OUT.t13 28.5655
R384 OUT.n4 OUT.t1 28.5655
R385 OUT.n0 OUT.t0 28.5655
R386 OUT.n0 OUT.t10 28.5655
R387 OUT.n18 OUT.t19 17.4005
R388 OUT.n18 OUT.t15 17.4005
R389 OUT.t8 OUT.n15 17.4005
R390 OUT.n15 OUT.t22 17.4005
R391 OUT.n14 OUT.n13 9.55736
R392 OUT OUT.n2 9.51046
R393 OUT OUT.n24 9.15531
R394 OUT OUT.n21 8.34995
R395 OUT.n10 OUT.n9 3.9555
R396 OUT.n6 OUT.n5 3.9555
R397 OUT.n23 OUT.n22 3.9555
R398 OUT OUT.n25 2.70196
R399 OUT.n21 OUT.n20 2.06216
R400 OUT.n21 OUT.n17 2.04399
R401 OUT.n24 OUT.n23 0.764437
R402 OUT.n20 OUT.n19 0.641024
R403 OUT.n17 OUT.n16 0.641024
R404 OUT.n14 OUT.n10 0.64003
R405 OUT.n5 OUT.n3 0.63421
R406 OUT.n6 OUT 0.62123
R407 OUT.n9 OUT.n7 0.617796
R408 OUT.n13 OUT.n11 0.61309
R409 OUT.n2 OUT.n1 0.594104
R410 OUT.n24 OUT.n14 0.474773
R411 OUT.n10 OUT.n6 0.355226
R412 OUT.n23 OUT 0.10188
R413 VIP.t2 VIP.t3 481.337
R414 VIP.n0 VIP.t1 240.865
R415 VIP VIP.t0 240.45
R416 VIP.t1 VIP.t2 237.144
R417 VIP.n2 VIP.n1 7.43383
R418 VIP.n2 VIP.n0 1.96558
R419 VIP VIP.n2 0.0594623
R420 VIP.n0 VIP 0.03175
R421 RS.n0 RS.t1 43.1877
R422 RS RS.t0 42.7848
R423 RS.n2 RS.n0 2.66873
R424 RS.n2 RS.n1 0.502858
R425 RS.n0 RS 0.234196
R426 RS RS.n2 0.00277273
R427 VIN.t2 VIN.t3 490.462
R428 VIN VIN.t0 245.508
R429 VIN.n0 VIN.t1 240.349
R430 VIN.t1 VIN.t2 237.144
R431 VIN.n2 VIN.n0 6.06934
R432 VIN.n0 VIN 4.59552
R433 VIN.n2 VIN.n1 0.50329
R434 VIN VIN.n2 0.00220455
C0 pmosdif_0.D5 pmosdif_0.D6 1.10858f
C1 pmosdif_0.D5 VIN 0.376877f
C2 pmosdif_0.D5 OUT 1.43031f
C3 pmoscs_0.D1 pmosdif_0.D5 1.46314f
C4 pmoscs_0.D2 VDD 4.12279f
C5 VIP VDD 0.856303f
C6 RS pmosdif_0.D5 0.033296f
C7 VIP pmosdif_0.D6 0.155604f
C8 VIP VIN 1.45283f
C9 OUT pmoscs_0.D2 0.065167f
C10 VIP OUT 0.669824f
C11 pmoscs_0.D1 pmoscs_0.D2 1.9701f
C12 VIP pmoscs_0.D1 0.01404f
C13 RS pmoscs_0.D2 0.66725f
C14 VIP RS 0.223097f
C15 pmosdif_0.D5 pmoscs_0.D2 1.70721f
C16 VIP pmosdif_0.D5 0.268208f
C17 pmosdif_0.D6 VDD 1.34306f
C18 VDD VIN 0.769669f
C19 OUT VDD 1.78349f
C20 pmosdif_0.D6 VIN 0.767919f
C21 OUT pmosdif_0.D6 2.76222f
C22 pmoscs_0.D1 VDD 1.3857f
C23 OUT VIN 0.156482f
C24 pmoscs_0.D1 pmosdif_0.D6 0.030356f
C25 RS VDD 0.278313f
C26 VIP pmoscs_0.D2 0.030428f
C27 pmoscs_0.D1 VIN 0.041257f
C28 RS pmosdif_0.D6 0.054178f
C29 pmoscs_0.D1 OUT 0.138692f
C30 RS VIN 0.046593f
C31 RS OUT 0.02749f
C32 pmosdif_0.D5 VDD 1.67295f
C33 RS pmoscs_0.D1 0.332322f
C34 VIN GND 0.875077f
C35 VIP GND 0.570435f
C36 OUT GND 4.105749f
C37 RS GND 1.40036f
C38 VDD GND 21.771132f
C39 pmosdif_0.D6 GND 6.930349f
C40 pmoscs_0.D1 GND 4.35654f
C41 pmoscs_0.D2 GND 3.113255f
C42 pmosdif_0.D5 GND 1.82057f
C43 OUT.n0 GND 0.013119f
C44 OUT.t11 GND 0.02334f
C45 OUT.t9 GND 0.01704f
C46 OUT.n1 GND 0.031436f
C47 OUT.n2 GND 0.177567f
C48 OUT.t12 GND 0.017238f
C49 OUT.n3 GND 0.03647f
C50 OUT.t13 GND 0.029711f
C51 OUT.n4 GND 0.013119f
C52 OUT.n5 GND 0.091486f
C53 OUT.n6 GND 0.107342f
C54 OUT.t5 GND 0.017061f
C55 OUT.n7 GND 0.031846f
C56 OUT.t6 GND 0.029716f
C57 OUT.n8 GND 0.013119f
C58 OUT.n9 GND 0.091504f
C59 OUT.n10 GND 0.108934f
C60 OUT.t4 GND 0.023334f
C61 OUT.t2 GND 0.017196f
C62 OUT.n11 GND 0.03594f
C63 OUT.n12 GND 0.013119f
C64 OUT.n13 GND 0.16969f
C65 OUT.n14 GND 0.120671f
C66 OUT.n15 GND 0.013847f
C67 OUT.t8 GND 0.028464f
C68 OUT.t7 GND 0.017037f
C69 OUT.n16 GND 0.036045f
C70 OUT.n17 GND 0.121732f
C71 OUT.n18 GND 0.013847f
C72 OUT.t16 GND 0.022086f
C73 OUT.t14 GND 0.016865f
C74 OUT.n19 GND 0.036152f
C75 OUT.n20 GND 0.120873f
C76 OUT.n21 GND 0.101674f
C77 OUT.t21 GND 0.022418f
C78 OUT.t20 GND 0.022418f
C79 OUT.n22 GND 0.118089f
C80 OUT.n23 GND 0.111872f
C81 OUT.n24 GND 0.275946f
C82 OUT.n25 GND 0.057442f
C83 pmosdif_0.D6.n0 GND 0.142102f
C84 pmosdif_0.D6.t29 GND 0.091392f
C85 pmosdif_0.D6.n1 GND 0.074296f
C86 pmosdif_0.D6.t30 GND 0.091422f
C87 pmosdif_0.D6.t10 GND 0.091423f
C88 pmosdif_0.D6.t16 GND 0.017428f
C89 pmosdif_0.D6.t14 GND 0.013444f
C90 pmosdif_0.D6.n2 GND 0.028441f
C91 pmosdif_0.D6.n3 GND 0.010927f
C92 pmosdif_0.D6.t25 GND 0.013444f
C93 pmosdif_0.D6.n4 GND 0.028441f
C94 pmosdif_0.D6.n5 GND 0.010352f
C95 pmosdif_0.D6.t13 GND 0.023446f
C96 pmosdif_0.D6.t12 GND 0.01357f
C97 pmosdif_0.D6.n6 GND 0.02836f
C98 pmosdif_0.D6.n7 GND 0.078432f
C99 pmosdif_0.D6.t21 GND 0.018411f
C100 pmosdif_0.D6.t19 GND 0.013641f
C101 pmosdif_0.D6.n8 GND 0.028774f
C102 pmosdif_0.D6.n9 GND 0.010352f
C103 pmosdif_0.D6.n10 GND 0.063307f
C104 pmosdif_0.D6.n11 GND 0.062589f
C105 pmosdif_0.D6.t24 GND 0.018411f
C106 pmosdif_0.D6.t22 GND 0.013588f
C107 pmosdif_0.D6.n12 GND 0.028678f
C108 pmosdif_0.D6.n13 GND 0.010352f
C109 pmosdif_0.D6.n14 GND 0.063314f
C110 pmosdif_0.D6.n15 GND 0.03893f
C111 pmosdif_0.D6.t17 GND 0.01357f
C112 pmosdif_0.D6.n16 GND 0.02836f
C113 pmosdif_0.D6.t18 GND 0.023446f
C114 pmosdif_0.D6.n17 GND 0.010352f
C115 pmosdif_0.D6.n18 GND 0.095015f
C116 pmosdif_0.D6.n19 GND 0.111006f
C117 pmosdif_0.D6.t27 GND 0.091422f
C118 pmosdif_0.D6.t4 GND 0.091423f
C119 pmosdif_0.D6.t9 GND 0.017676f
C120 pmosdif_0.D6.t7 GND 0.017676f
C121 pmosdif_0.D6.n20 GND 0.077997f
C122 pmosdif_0.D6.t8 GND 0.090922f
C123 pmosdif_0.D6.t6 GND 0.090882f
C124 pmosdif_0.D6.n21 GND 0.07812f
C125 pmosdif_0.D6.n22 GND 0.021392f
C126 pmosdif_0.D6.t28 GND 0.091392f
C127 pmosdif_0.D6.n23 GND 0.074296f
C128 pmosdif_0.D6.n24 GND 0.132956f
C129 pmosdif_0.D6.n25 GND 0.045534f
C130 pmosdif_0.D6.t26 GND 0.022461f
C131 pmosdif_0.D6.n26 GND 0.010927f
C132 pmosdif_0.D6.n27 GND 0.13972f
C133 pmoscs_0.D2.n0 GND 0.355946f
C134 pmoscs_0.D2.n1 GND 0.311868f
C135 pmoscs_0.D2.t1 GND 0.042352f
C136 pmoscs_0.D2.t0 GND 0.024868f
C137 pmoscs_0.D2.n2 GND 0.06592f
C138 pmoscs_0.D2.t2 GND 0.04276f
C139 pmoscs_0.D2.t16 GND 0.042794f
C140 pmoscs_0.D2.t15 GND 0.042794f
C141 pmoscs_0.D2.t8 GND 0.041073f
C142 pmoscs_0.D2.n3 GND 0.031752f
C143 pmoscs_0.D2.t9 GND 0.0247f
C144 pmoscs_0.D2.n4 GND 0.029288f
C145 pmoscs_0.D2.t11 GND 0.151815f
C146 pmoscs_0.D2.n5 GND 0.041317f
C147 pmoscs_0.D2.t5 GND 0.045069f
C148 pmoscs_0.D2.t3 GND 0.025115f
C149 pmoscs_0.D2.n6 GND 0.070683f
C150 pmoscs_0.D2.t14 GND 0.012298f
C151 pmoscs_0.D2.t4 GND 0.012298f
C152 pmoscs_0.D2.n7 GND 0.025411f
C153 pmoscs_0.D2.n8 GND 0.192307f
C154 pmoscs_0.D2.n9 GND 0.108634f
C155 pmoscs_0.D2.t17 GND 0.274453f
C156 pmoscs_0.D2.t18 GND 0.22186f
C157 pmoscs_0.D2.t13 GND 0.182496f
C158 pmoscs_0.D2.n10 GND 0.076574f
C159 pmoscs_0.D2.n11 GND 0.09803f
C160 pmoscs_0.D2.t20 GND 0.274453f
C161 pmoscs_0.D2.t19 GND 0.221647f
C162 pmoscs_0.D2.n12 GND 0.098031f
C163 pmoscs_0.D2.n13 GND 0.076682f
C164 pmoscs_0.D2.t10 GND 0.056777f
C165 pmoscs_0.D2.t12 GND 0.012298f
C166 pmoscs_0.D2.n14 GND 0.025411f
C167 pmoscs_0.D2.n15 GND 0.17988f
C168 pmoscs_0.D2.n16 GND 0.088162f
C169 pmoscs_0.D2.t6 GND 0.024459f
C170 pmoscs_0.D2.n17 GND 0.026596f
C171 pmoscs_0.D2.n18 GND 0.017652f
C172 pmoscs_0.D2.t7 GND 0.04276f
C173 VDD.n0 GND 0.015139f
C174 VDD.n1 GND 0.02902f
C175 VDD.n2 GND 0.02902f
C176 VDD.n3 GND 0.02902f
C177 VDD.t3 GND 0.184884f
C178 VDD.n4 GND 0.028663f
C179 VDD.n5 GND 0.184914f
C180 VDD.t2 GND 0.199096f
C181 VDD.t5 GND 0.139522f
C182 VDD.n6 GND 0.055671f
C183 VDD.t0 GND 0.137461f
C184 VDD.n7 GND 0.280939f
C185 VDD.n8 GND 0.174906f
C186 VDD.n9 GND 0.028674f
C187 VDD.n10 GND 0.028061f
C188 VDD.n11 GND 0.014638f
C189 VDD.n12 GND 0.030591f
C190 VDD.n13 GND 0.030605f
C191 VDD.n14 GND 0.212517f
C192 VDD.n15 GND 0.033895f
C193 VDD.t4 GND 0.266823f
C194 VDD.t6 GND 0.236491f
C195 VDD.t16 GND 0.057404f
C196 VDD.n16 GND 0.018348f
C197 VDD.t19 GND 0.014676f
C198 VDD.n22 GND 0.033325f
C199 VDD.t14 GND 0.057404f
C200 VDD.n23 GND 0.018648f
C201 VDD.n24 GND 0.025935f
C202 VDD.n26 GND 0.021353f
C203 VDD.n28 GND 0.021365f
C204 VDD.n29 GND 0.025827f
C205 VDD.n32 GND 0.032988f
C206 VDD.t22 GND 0.011497f
C207 VDD.n36 GND 0.017194f
C208 VDD.n37 GND 0.020318f
C209 VDD.n38 GND 0.034188f
C210 VDD.n39 GND 0.199274f
C211 VDD.t1 GND 0.249062f
C212 VDD.t8 GND 0.236491f
C213 VDD.n40 GND 0.193654f
C214 VDD.n41 GND 0.102139f
C215 VDD.n42 GND 0.034207f
C216 VDD.n43 GND 0.020314f
C217 VDD.n44 GND 0.017178f
C218 VDD.n45 GND 0.028214f
C219 VDD.n46 GND 0.044476f
C220 VDD.n47 GND 0.018517f
.ends

