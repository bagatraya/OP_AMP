magic
tech sky130A
magscale 1 2
timestamp 1729219841
<< psubdiff >>
rect -176 518 -111 552
rect 1390 518 1450 552
rect -176 492 -142 518
rect 1416 492 1450 518
rect -176 -614 -142 -588
rect 1416 -614 1450 -588
rect -176 -648 -111 -614
rect 1390 -648 1450 -614
<< psubdiffcont >>
rect -111 518 1390 552
rect -176 -588 -142 492
rect 1416 -588 1450 492
rect -111 -648 1390 -614
<< poly >>
rect -30 66 0 88
rect -92 50 0 66
rect -92 16 -76 50
rect -42 16 0 50
rect -92 0 0 16
rect 1272 66 1302 88
rect 1272 50 1364 66
rect 1272 16 1314 50
rect 1348 16 1364 50
rect 1272 0 1364 16
rect -30 -1 0 0
rect -92 -112 0 -96
rect -92 -146 -76 -112
rect -42 -146 0 -112
rect -92 -162 0 -146
rect -30 -184 0 -162
rect 1272 -112 1364 -96
rect 1272 -146 1314 -112
rect 1348 -146 1364 -112
rect 1272 -162 1364 -146
rect 1272 -184 1302 -162
<< polycont >>
rect -76 16 -42 50
rect 1314 16 1348 50
rect -76 -146 -42 -112
rect 1314 -146 1348 -112
<< locali >>
rect -176 518 -111 552
rect 1390 518 1450 552
rect -176 492 -142 518
rect 1416 492 1450 518
rect -76 50 -42 100
rect 1314 50 1348 100
rect -92 16 -76 50
rect -42 16 -26 50
rect 1298 16 1314 50
rect 1348 16 1364 50
rect -92 -146 -76 -112
rect -42 -146 -26 -112
rect 1298 -146 1314 -112
rect 1348 -146 1364 -112
rect -76 -186 -42 -146
rect 1314 -196 1348 -146
rect -176 -614 -142 -588
rect 1416 -614 1450 -588
rect -176 -648 -111 -614
rect 1390 -648 1450 -614
<< viali >>
rect -76 16 -42 50
rect 1314 16 1348 50
rect -76 -146 -42 -112
rect 1314 -146 1348 -112
rect 277 -614 330 -613
rect 941 -614 994 -613
rect 277 -648 330 -614
rect 941 -648 994 -614
<< metal1 >>
rect 591 455 601 466
rect -39 407 601 455
rect -39 288 9 407
rect 591 396 601 407
rect 671 455 681 466
rect 1064 455 1312 456
rect 671 407 1312 455
rect 671 396 681 407
rect 1263 288 1312 407
rect -82 88 52 288
rect 224 88 384 288
rect -76 56 -42 88
rect -88 50 -30 56
rect -88 16 -76 50
rect -42 16 -30 50
rect -88 10 -30 16
rect 64 7 74 59
rect 202 7 212 59
rect -88 -112 -30 -106
rect -88 -146 -76 -112
rect -42 -146 -30 -112
rect -88 -152 -30 -146
rect -76 -186 -42 -152
rect 64 -157 74 -105
rect 202 -157 212 -105
rect 280 -184 328 88
rect 556 86 716 286
rect 888 88 1048 288
rect 1220 88 1354 288
rect 612 57 660 86
rect 604 55 610 57
rect 470 7 610 55
rect 604 5 610 7
rect 662 55 668 57
rect 662 7 801 55
rect 662 5 668 7
rect 396 -155 406 -103
rect 534 -155 544 -103
rect 728 -155 738 -103
rect 866 -155 876 -103
rect 944 -184 992 88
rect 1060 7 1070 59
rect 1198 7 1208 59
rect 1314 56 1348 88
rect 1302 50 1360 56
rect 1302 16 1314 50
rect 1348 16 1360 50
rect 1302 10 1360 16
rect 1060 -157 1070 -105
rect 1198 -157 1208 -105
rect 1302 -112 1360 -106
rect 1302 -146 1314 -112
rect 1348 -146 1360 -112
rect 1302 -152 1360 -146
rect -82 -198 52 -186
rect -82 -374 -41 -198
rect 11 -374 52 -198
rect -82 -386 52 -374
rect 224 -196 384 -184
rect 224 -372 278 -196
rect 330 -372 384 -196
rect 224 -384 384 -372
rect 556 -196 716 -184
rect 556 -372 608 -196
rect 664 -372 716 -196
rect 556 -384 716 -372
rect 888 -196 1048 -184
rect 1314 -186 1348 -152
rect 888 -372 942 -196
rect 994 -372 1048 -196
rect 888 -384 1048 -372
rect 1220 -200 1354 -186
rect 1220 -367 1261 -200
rect 1313 -367 1354 -200
rect 1220 -386 1354 -367
rect -41 -510 11 -386
rect 1261 -510 1313 -386
rect -41 -562 1313 -510
rect 267 -607 277 -604
rect 265 -654 277 -607
rect 329 -607 339 -604
rect 932 -607 942 -604
rect 329 -613 342 -607
rect 330 -648 342 -613
rect 267 -656 277 -654
rect 329 -654 342 -648
rect 929 -613 942 -607
rect 994 -607 1004 -604
rect 929 -648 941 -613
rect 929 -654 942 -648
rect 329 -656 339 -654
rect 932 -656 942 -654
rect 994 -654 1006 -607
rect 994 -656 1004 -654
<< via1 >>
rect 601 396 671 466
rect 74 7 202 59
rect 74 -157 202 -105
rect 610 5 662 57
rect 406 -155 534 -103
rect 738 -155 866 -103
rect 1070 7 1198 59
rect 1070 -157 1198 -105
rect -41 -374 11 -198
rect 278 -372 330 -196
rect 608 -372 664 -196
rect 942 -372 994 -196
rect 1261 -367 1313 -200
rect 277 -613 329 -604
rect 277 -648 329 -613
rect 277 -656 329 -648
rect 942 -613 994 -604
rect 942 -648 994 -613
rect 942 -656 994 -648
<< metal2 >>
rect 601 466 671 476
rect 601 386 671 396
rect 74 59 202 69
rect 74 -22 202 7
rect 610 57 662 63
rect 610 -22 662 5
rect 1070 59 1198 69
rect 1070 -22 1198 7
rect -41 -74 1313 -22
rect -41 -198 11 -74
rect 74 -105 202 -74
rect 74 -167 202 -157
rect 406 -103 534 -74
rect 406 -165 534 -155
rect 738 -103 866 -74
rect 738 -165 866 -155
rect 1070 -105 1198 -74
rect 1070 -167 1198 -157
rect 278 -196 330 -186
rect -41 -382 11 -374
rect 277 -372 278 -348
rect 277 -382 330 -372
rect 608 -196 664 -186
rect 608 -382 664 -372
rect 942 -196 994 -186
rect 277 -509 329 -382
rect 942 -509 994 -372
rect 1261 -200 1313 -74
rect 1261 -378 1313 -367
rect 277 -561 994 -509
rect 277 -604 329 -561
rect 277 -666 329 -656
rect 942 -604 994 -561
rect 942 -666 994 -656
<< via2 >>
rect 606 401 666 461
rect 608 -372 664 -196
<< metal3 >>
rect 601 461 671 466
rect 601 401 606 461
rect 666 401 671 461
rect 601 396 671 401
rect 606 -191 666 396
rect 598 -196 674 -191
rect 598 -372 608 -196
rect 664 -372 674 -196
rect 598 -377 674 -372
use sky130_fd_pr__nfet_01v8_6H9P4D  sky130_fd_pr__nfet_01v8_6H9P4D_0
timestamp 1729213091
transform 1 0 -15 0 1 188
box -73 -126 73 126
use sky130_fd_pr__nfet_01v8_6H9P4D  sky130_fd_pr__nfet_01v8_6H9P4D_1
timestamp 1729213091
transform 1 0 -15 0 1 -284
box -73 -126 73 126
use sky130_fd_pr__nfet_01v8_6H9P4D  sky130_fd_pr__nfet_01v8_6H9P4D_2
timestamp 1729213091
transform 1 0 1287 0 1 188
box -73 -126 73 126
use sky130_fd_pr__nfet_01v8_6H9P4D  sky130_fd_pr__nfet_01v8_6H9P4D_3
timestamp 1729213091
transform 1 0 1287 0 1 -284
box -73 -126 73 126
use sky130_fd_pr__nfet_01v8_DB328X  sky130_fd_pr__nfet_01v8_DB328X_0
timestamp 1729208699
transform 1 0 636 0 1 188
box -636 -188 636 188
use sky130_fd_pr__nfet_01v8_DB328X  sky130_fd_pr__nfet_01v8_DB328X_1
timestamp 1729208699
transform 1 0 636 0 1 -284
box -636 -188 636 188
<< labels >>
flabel metal3 632 -135 632 -135 0 FreeSans 480 0 0 0 OUT
port 1 nsew
flabel metal2 135 -48 135 -48 0 FreeSans 480 0 0 0 D6
port 2 nsew
flabel metal2 968 -454 968 -454 0 FreeSans 480 0 0 0 GND
port 0 nsew
<< end >>
