magic
tech sky130A
magscale 1 2
timestamp 1729208699
<< nmos >>
rect -189 109 -29 309
rect 29 109 189 309
rect -189 -309 -29 -109
rect 29 -309 189 -109
<< ndiff >>
rect -247 297 -189 309
rect -247 121 -235 297
rect -201 121 -189 297
rect -247 109 -189 121
rect -29 297 29 309
rect -29 121 -17 297
rect 17 121 29 297
rect -29 109 29 121
rect 189 297 247 309
rect 189 121 201 297
rect 235 121 247 297
rect 189 109 247 121
rect -247 -121 -189 -109
rect -247 -297 -235 -121
rect -201 -297 -189 -121
rect -247 -309 -189 -297
rect -29 -121 29 -109
rect -29 -297 -17 -121
rect 17 -297 29 -121
rect -29 -309 29 -297
rect 189 -121 247 -109
rect 189 -297 201 -121
rect 235 -297 247 -121
rect 189 -309 247 -297
<< ndiffc >>
rect -235 121 -201 297
rect -17 121 17 297
rect 201 121 235 297
rect -235 -297 -201 -121
rect -17 -297 17 -121
rect 201 -297 235 -121
<< poly >>
rect -189 381 -29 397
rect -189 347 -173 381
rect -45 347 -29 381
rect -189 309 -29 347
rect 29 381 189 397
rect 29 347 45 381
rect 173 347 189 381
rect 29 309 189 347
rect -189 71 -29 109
rect -189 37 -173 71
rect -45 37 -29 71
rect -189 21 -29 37
rect 29 71 189 109
rect 29 37 45 71
rect 173 37 189 71
rect 29 21 189 37
rect -189 -37 -29 -21
rect -189 -71 -173 -37
rect -45 -71 -29 -37
rect -189 -109 -29 -71
rect 29 -37 189 -21
rect 29 -71 45 -37
rect 173 -71 189 -37
rect 29 -109 189 -71
rect -189 -347 -29 -309
rect -189 -381 -173 -347
rect -45 -381 -29 -347
rect -189 -397 -29 -381
rect 29 -347 189 -309
rect 29 -381 45 -347
rect 173 -381 189 -347
rect 29 -397 189 -381
<< polycont >>
rect -173 347 -45 381
rect 45 347 173 381
rect -173 37 -45 71
rect 45 37 173 71
rect -173 -71 -45 -37
rect 45 -71 173 -37
rect -173 -381 -45 -347
rect 45 -381 173 -347
<< locali >>
rect -189 347 -173 381
rect -45 347 -29 381
rect 29 347 45 381
rect 173 347 189 381
rect -235 297 -201 313
rect -235 105 -201 121
rect -17 297 17 313
rect -17 105 17 121
rect 201 297 235 313
rect 201 105 235 121
rect -189 37 -173 71
rect -45 37 -29 71
rect 29 37 45 71
rect 173 37 189 71
rect -189 -71 -173 -37
rect -45 -71 -29 -37
rect 29 -71 45 -37
rect 173 -71 189 -37
rect -235 -121 -201 -105
rect -235 -313 -201 -297
rect -17 -121 17 -105
rect -17 -313 17 -297
rect 201 -121 235 -105
rect 201 -313 235 -297
rect -189 -381 -173 -347
rect -45 -381 -29 -347
rect 29 -381 45 -347
rect 173 -381 189 -347
<< viali >>
rect -173 347 -45 381
rect 45 347 173 381
rect -235 121 -201 297
rect -17 121 17 297
rect 201 121 235 297
rect -173 37 -45 71
rect 45 37 173 71
rect -173 -71 -45 -37
rect 45 -71 173 -37
rect -235 -297 -201 -121
rect -17 -297 17 -121
rect 201 -297 235 -121
rect -173 -381 -45 -347
rect 45 -381 173 -347
<< metal1 >>
rect -185 381 -33 387
rect -185 347 -173 381
rect -45 347 -33 381
rect -185 341 -33 347
rect 33 381 185 387
rect 33 347 45 381
rect 173 347 185 381
rect 33 341 185 347
rect -241 297 -195 309
rect -241 121 -235 297
rect -201 121 -195 297
rect -241 109 -195 121
rect -23 297 23 309
rect -23 121 -17 297
rect 17 121 23 297
rect -23 109 23 121
rect 195 297 241 309
rect 195 121 201 297
rect 235 121 241 297
rect 195 109 241 121
rect -185 71 -33 77
rect -185 37 -173 71
rect -45 37 -33 71
rect -185 31 -33 37
rect 33 71 185 77
rect 33 37 45 71
rect 173 37 185 71
rect 33 31 185 37
rect -185 -37 -33 -31
rect -185 -71 -173 -37
rect -45 -71 -33 -37
rect -185 -77 -33 -71
rect 33 -37 185 -31
rect 33 -71 45 -37
rect 173 -71 185 -37
rect 33 -77 185 -71
rect -241 -121 -195 -109
rect -241 -297 -235 -121
rect -201 -297 -195 -121
rect -241 -309 -195 -297
rect -23 -121 23 -109
rect -23 -297 -17 -121
rect 17 -297 23 -121
rect -23 -309 23 -297
rect 195 -121 241 -109
rect 195 -297 201 -121
rect 235 -297 241 -121
rect 195 -309 241 -297
rect -185 -347 -33 -341
rect -185 -381 -173 -347
rect -45 -381 -33 -347
rect -185 -387 -33 -381
rect 33 -347 185 -341
rect 33 -381 45 -347
rect 173 -381 185 -347
rect 33 -387 185 -381
<< properties >>
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 1 l 0.8 m 2 nf 2 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
