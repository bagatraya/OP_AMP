magic
tech sky130A
magscale 1 2
timestamp 1729236107
<< nwell >>
rect -323 2866 678 3039
rect 2418 2469 3224 3040
<< viali >>
rect 2131 2612 2331 2812
rect 2130 2355 2330 2555
rect 2127 2085 2327 2285
rect 2125 1807 2325 2007
rect 1977 1617 2012 1679
rect 2125 1537 2325 1737
rect 2125 1271 2325 1471
rect 1402 1202 1448 1239
<< metal1 >>
rect 498 2866 2706 2922
rect 498 2798 554 2866
rect 2201 2818 2257 2866
rect 2119 2812 2343 2818
rect 2119 2612 2131 2812
rect 2331 2612 2343 2812
rect 2119 2606 2343 2612
rect 2118 2555 2342 2561
rect 2118 2355 2130 2555
rect 2330 2355 2342 2555
rect 2650 2470 2706 2866
rect 2118 2349 2342 2355
rect 2115 2285 2339 2291
rect 642 2169 652 2248
rect 726 2241 736 2248
rect 726 2178 868 2241
rect 726 2169 736 2178
rect 2115 2085 2127 2285
rect 2327 2215 2339 2285
rect 2327 2163 2450 2215
rect 2327 2085 2339 2163
rect 2115 2079 2339 2085
rect 368 2028 884 2066
rect 2113 2007 2337 2013
rect 2113 1807 2125 2007
rect 2325 1807 2337 2007
rect 2113 1801 2337 1807
rect 2398 1781 2450 2163
rect 2113 1737 2337 1743
rect 1971 1679 2018 1691
rect 2113 1679 2125 1737
rect 1971 1617 1977 1679
rect 2012 1617 2125 1679
rect 1971 1615 2125 1617
rect 1971 1605 2018 1615
rect 2113 1537 2125 1615
rect 2325 1537 2337 1737
rect 2398 1729 2773 1781
rect 2393 1646 2399 1698
rect 2451 1646 2797 1698
rect 2113 1531 2337 1537
rect 2113 1471 2337 1477
rect 1402 1245 1450 1458
rect 2113 1271 2125 1471
rect 2325 1404 2337 1471
rect 2325 1338 2436 1404
rect 2325 1271 2337 1338
rect 2113 1265 2337 1271
rect 1390 1239 1460 1245
rect 1390 1202 1402 1239
rect 1448 1202 1460 1239
rect 1390 1196 1460 1202
rect 2370 1156 2436 1338
rect 2363 1090 2373 1156
rect 2439 1090 2449 1156
<< via1 >>
rect 2130 2355 2330 2555
rect 652 2169 726 2248
rect 2125 1807 2325 2007
rect 2399 1646 2451 1698
rect 2373 1090 2439 1156
<< metal2 >>
rect 2130 2555 2330 2565
rect 2035 2435 2130 2481
rect 652 2248 726 2258
rect 652 2159 726 2169
rect 2035 2156 2081 2435
rect 2130 2345 2330 2355
rect 1402 2110 2081 2156
rect 2125 2007 2325 2017
rect 2325 1879 2451 1931
rect 2125 1797 2325 1807
rect 2399 1698 2451 1879
rect 2721 1739 2772 1772
rect 2399 1640 2451 1646
rect 887 1368 980 1378
rect 507 1295 887 1356
rect 887 1276 980 1286
rect 2373 1156 2439 1166
rect 2369 1095 2373 1151
rect 2439 1095 2443 1151
rect 2373 1080 2439 1090
rect 2167 610 2603 662
<< via2 >>
rect 652 2169 726 2248
rect 887 1286 980 1368
rect 2373 1090 2439 1156
<< metal3 >>
rect 642 2248 736 2253
rect 642 2169 652 2248
rect 726 2169 736 2248
rect 642 2164 736 2169
rect 660 1467 723 2164
rect 413 1404 723 1467
rect 877 1368 990 1373
rect 877 1286 887 1368
rect 980 1355 990 1368
rect 980 1294 2856 1355
rect 980 1286 990 1294
rect 877 1281 990 1286
rect 2363 1156 2449 1161
rect 2363 1090 2373 1156
rect 2439 1090 2449 1156
rect 2363 1085 2449 1090
rect 1508 180 1574 312
rect 2373 180 2439 1085
rect 1508 114 3044 180
use nmoscs  nmoscs_0
timestamp 1729179123
transform 1 0 1024 0 1 2233
box -290 -815 988 605
use nmosdif  nmosdif_0
timestamp 1729219841
transform 1 0 906 0 1 684
box -176 -666 1450 552
use pmoscs  pmoscs_0
timestamp 1729157559
transform 1 0 -353 0 1 480
box 34 -480 1032 2387
use pmosdif  pmosdif_0
timestamp 1729197635
transform 1 0 2101 0 1 1610
box 324 -1596 1124 912
<< labels >>
flabel viali 2232 1397 2234 1398 0 FreeSans 800 0 0 0 OUT
port 0 nsew
flabel viali 2221 1640 2223 1641 0 FreeSans 800 0 0 0 GND
port 1 nsew
flabel via1 2222 1912 2222 1912 0 FreeSans 800 0 0 0 VIN
port 2 nsew
flabel viali 2127 2085 2327 2285 0 FreeSans 800 0 0 0 VIP
port 3 nsew
flabel via1 2234 2458 2234 2458 0 FreeSans 800 0 0 0 RS
port 4 nsew
flabel viali 2224 2716 2224 2716 0 FreeSans 800 0 0 0 VDD
port 6 nsew
<< end >>
