magic
tech sky130A
magscale 1 2
timestamp 1729189057
<< nwell >>
rect -223 -200 223 200
<< pmos >>
rect -129 -100 -29 100
rect 29 -100 129 100
<< pdiff >>
rect -187 88 -129 100
rect -187 -88 -175 88
rect -141 -88 -129 88
rect -187 -100 -129 -88
rect -29 88 29 100
rect -29 -88 -17 88
rect 17 -88 29 88
rect -29 -100 29 -88
rect 129 88 187 100
rect 129 -88 141 88
rect 175 -88 187 88
rect 129 -100 187 -88
<< pdiffc >>
rect -175 -88 -141 88
rect -17 -88 17 88
rect 141 -88 175 88
<< poly >>
rect -126 181 -32 197
rect -126 164 -110 181
rect -129 147 -110 164
rect -48 164 -32 181
rect 32 181 126 197
rect 32 164 48 181
rect -48 147 -29 164
rect -129 100 -29 147
rect 29 147 48 164
rect 110 164 126 181
rect 110 147 129 164
rect 29 100 129 147
rect -129 -147 -29 -100
rect -129 -164 -110 -147
rect -126 -181 -110 -164
rect -48 -164 -29 -147
rect 29 -147 129 -100
rect 29 -164 48 -147
rect -48 -181 -32 -164
rect -126 -197 -32 -181
rect 32 -181 48 -164
rect 110 -164 129 -147
rect 110 -181 126 -164
rect 32 -197 126 -181
<< polycont >>
rect -110 147 -48 181
rect 48 147 110 181
rect -110 -181 -48 -147
rect 48 -181 110 -147
<< locali >>
rect -126 147 -110 181
rect -48 147 -32 181
rect 32 147 48 181
rect 110 147 126 181
rect -175 88 -141 104
rect -175 -104 -141 -88
rect -17 88 17 104
rect -17 -104 17 -88
rect 141 88 175 104
rect 141 -104 175 -88
rect -126 -181 -110 -147
rect -48 -181 -32 -147
rect 32 -181 48 -147
rect 110 -181 126 -147
<< viali >>
rect -106 147 -52 181
rect 52 147 106 181
rect -175 -88 -141 88
rect -17 -88 17 88
rect 141 -88 175 88
rect -106 -181 -52 -147
rect 52 -181 106 -147
<< metal1 >>
rect -118 181 -40 187
rect -118 147 -106 181
rect -52 147 -40 181
rect -118 141 -40 147
rect 40 181 118 187
rect 40 147 52 181
rect 106 147 118 181
rect 40 141 118 147
rect -181 88 -135 100
rect -181 -88 -175 88
rect -141 -88 -135 88
rect -181 -100 -135 -88
rect -23 88 23 100
rect -23 -88 -17 88
rect 17 -88 23 88
rect -23 -100 23 -88
rect 135 88 181 100
rect 135 -88 141 88
rect 175 -88 181 88
rect 135 -100 181 -88
rect -118 -147 -40 -141
rect -118 -181 -106 -147
rect -52 -181 -40 -147
rect -118 -187 -40 -181
rect 40 -147 118 -141
rect 40 -181 52 -147
rect 106 -181 118 -147
rect 40 -187 118 -181
<< properties >>
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 1 l 0.5 m 1 nf 2 diffcov 100 polycov 90 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 80 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
