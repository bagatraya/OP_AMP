magic
tech sky130A
magscale 1 2
timestamp 1729157559
<< nwell >>
rect 34 -480 1032 2387
<< nsubdiff >>
rect 70 2317 132 2351
rect 936 2317 996 2351
rect 70 2289 104 2317
rect 962 2289 996 2317
rect 70 -410 104 -382
rect 962 -410 996 -382
rect 70 -444 132 -410
rect 936 -444 996 -410
<< nsubdiffcont >>
rect 132 2317 936 2351
rect 70 -382 104 2289
rect 962 -382 996 2289
rect 132 -444 936 -410
<< poly >>
rect 154 2277 246 2293
rect 154 2243 170 2277
rect 204 2243 246 2277
rect 154 2227 246 2243
rect 216 2196 246 2227
rect 820 2277 912 2293
rect 820 2243 862 2277
rect 896 2243 912 2277
rect 820 2227 912 2243
rect 820 2196 850 2227
rect 304 1598 504 1699
rect 154 1582 246 1598
rect 154 1548 170 1582
rect 204 1548 246 1582
rect 154 1532 246 1548
rect 216 1501 246 1532
rect 820 1583 912 1599
rect 820 1549 862 1583
rect 896 1549 912 1583
rect 820 1533 912 1549
rect 820 1502 850 1533
rect 304 903 762 1004
rect 216 375 246 406
rect 154 359 246 375
rect 154 325 170 359
rect 204 325 246 359
rect 154 309 246 325
rect 820 375 850 406
rect 820 359 912 375
rect 820 325 862 359
rect 896 325 912 359
rect 820 309 912 325
rect 562 208 762 309
rect 216 -320 246 -278
rect 154 -336 246 -320
rect 154 -370 170 -336
rect 204 -370 246 -336
rect 154 -385 246 -370
rect 820 -320 850 -289
rect 820 -336 912 -320
rect 820 -370 862 -336
rect 896 -370 912 -336
rect 820 -385 912 -370
rect 846 -386 912 -385
<< polycont >>
rect 170 2243 204 2277
rect 862 2243 896 2277
rect 170 1548 204 1582
rect 862 1549 896 1583
rect 170 325 204 359
rect 862 325 896 359
rect 170 -370 204 -336
rect 862 -370 896 -336
<< locali >>
rect 70 2317 132 2351
rect 936 2317 996 2351
rect 70 2289 104 2317
rect 962 2289 996 2317
rect 154 2243 170 2277
rect 204 2243 220 2277
rect 846 2243 862 2277
rect 896 2243 912 2277
rect 170 2196 204 2243
rect 862 2200 896 2243
rect 158 1796 218 2196
rect 154 1548 170 1582
rect 204 1548 220 1582
rect 846 1549 862 1583
rect 896 1549 912 1583
rect 170 1502 204 1548
rect 862 1502 896 1549
rect 160 1102 212 1502
rect 246 1102 306 1502
rect 766 1102 818 1502
rect 854 1102 906 1502
rect 160 408 212 808
rect 250 408 302 808
rect 768 408 820 808
rect 170 359 204 408
rect 862 359 896 418
rect 154 325 170 359
rect 204 325 220 359
rect 846 325 862 359
rect 896 325 912 359
rect 170 -336 204 -277
rect 850 -288 902 112
rect 862 -336 896 -288
rect 154 -370 170 -336
rect 204 -370 220 -336
rect 846 -370 862 -336
rect 896 -370 912 -336
rect 70 -410 104 -382
rect 962 -410 996 -382
rect 70 -444 132 -410
rect 936 -444 996 -410
<< viali >>
rect 861 2351 896 2352
rect 861 2317 896 2351
rect 170 2243 204 2277
rect 862 2243 896 2277
rect 170 1548 204 1582
rect 862 1549 896 1583
rect 170 325 204 359
rect 862 325 896 359
rect 170 -370 204 -336
rect 862 -370 896 -336
rect 170 -444 204 -410
<< metal1 >>
rect 849 2352 908 2358
rect 849 2317 861 2352
rect 896 2317 908 2352
rect 849 2311 908 2317
rect 862 2283 896 2311
rect 158 2277 216 2283
rect 158 2243 170 2277
rect 204 2243 216 2277
rect 158 2237 216 2243
rect 850 2277 908 2283
rect 850 2243 862 2277
rect 896 2243 908 2277
rect 850 2237 908 2243
rect 170 2198 204 2237
rect 165 2197 216 2198
rect 158 2185 304 2197
rect 151 1809 161 2185
rect 213 1809 304 2185
rect 158 1797 304 1809
rect 510 1756 556 2198
rect 862 2196 896 2237
rect 768 1796 902 2196
rect 768 1756 816 1796
rect 510 1708 816 1756
rect 158 1582 216 1588
rect 158 1548 170 1582
rect 204 1548 216 1582
rect 158 1542 216 1548
rect 170 1501 204 1542
rect 159 1488 306 1500
rect 159 1112 248 1488
rect 300 1112 310 1488
rect 159 1102 306 1112
rect 243 844 249 896
rect 301 844 475 896
rect 158 794 305 808
rect 158 418 249 794
rect 301 418 305 794
rect 158 407 305 418
rect 163 406 215 407
rect 248 406 304 407
rect 164 365 215 406
rect 158 359 216 365
rect 158 325 170 359
rect 204 325 216 359
rect 158 319 216 325
rect 510 198 556 1708
rect 850 1583 908 1589
rect 850 1549 862 1583
rect 896 1549 908 1583
rect 850 1543 908 1549
rect 862 1502 896 1543
rect 762 1501 908 1502
rect 756 1489 908 1501
rect 755 1113 765 1489
rect 817 1113 908 1489
rect 756 1101 908 1113
rect 765 1063 817 1069
rect 591 1011 765 1063
rect 765 1005 817 1011
rect 850 806 901 807
rect 761 794 908 806
rect 754 418 764 794
rect 816 418 908 794
rect 761 407 908 418
rect 850 406 904 407
rect 851 365 904 406
rect 850 359 908 365
rect 850 325 862 359
rect 896 325 908 359
rect 850 319 908 325
rect 252 152 556 198
rect 252 111 298 152
rect 164 -289 298 111
rect 510 -289 556 152
rect 853 111 901 115
rect 762 100 908 111
rect 762 -276 853 100
rect 905 -276 915 100
rect 762 -289 908 -276
rect 164 -330 210 -289
rect 853 -330 901 -289
rect 158 -336 216 -330
rect 158 -370 170 -336
rect 204 -370 216 -336
rect 158 -376 216 -370
rect 850 -336 908 -330
rect 850 -370 862 -336
rect 896 -370 908 -336
rect 850 -376 908 -370
rect 165 -404 210 -376
rect 158 -410 216 -404
rect 158 -444 170 -410
rect 204 -444 216 -410
rect 158 -450 216 -444
<< via1 >>
rect 161 1809 213 2185
rect 248 1112 300 1488
rect 249 844 301 896
rect 249 418 301 794
rect 765 1113 817 1489
rect 765 1011 817 1063
rect 764 418 816 794
rect 853 -276 905 100
<< metal2 >>
rect 161 2185 213 2195
rect 161 1687 213 1809
rect 159 1677 215 1687
rect 159 1611 215 1621
rect 849 1679 909 1688
rect 160 298 212 1611
rect 849 1610 909 1619
rect 247 1489 303 1499
rect 247 1112 248 1113
rect 300 1112 303 1113
rect 247 1103 303 1112
rect 765 1489 817 1499
rect 248 1102 300 1103
rect 765 1063 817 1113
rect 759 1011 765 1063
rect 817 1011 823 1063
rect 765 981 817 1011
rect 249 929 817 981
rect 249 896 301 929
rect 249 794 301 844
rect 768 807 825 817
rect 249 408 301 418
rect 764 794 768 804
rect 764 408 768 418
rect 768 396 825 406
rect 157 289 217 298
rect 853 297 905 1610
rect 157 220 217 229
rect 851 287 907 297
rect 851 221 907 231
rect 853 100 905 221
rect 853 -284 905 -276
<< via2 >>
rect 159 1621 215 1677
rect 849 1619 909 1679
rect 247 1488 303 1489
rect 247 1113 248 1488
rect 248 1113 300 1488
rect 300 1113 303 1488
rect 768 794 825 807
rect 768 418 816 794
rect 816 418 825 794
rect 768 406 825 418
rect 157 229 217 289
rect 851 231 907 287
<< metal3 >>
rect 149 1679 225 1682
rect 844 1679 914 1684
rect 149 1677 849 1679
rect 149 1621 159 1677
rect 215 1621 849 1677
rect 149 1619 849 1621
rect 909 1619 914 1679
rect 149 1616 225 1619
rect 844 1614 914 1619
rect 237 1489 313 1494
rect 237 1113 247 1489
rect 303 1113 313 1489
rect 237 1108 313 1113
rect 243 987 306 1108
rect 243 924 829 987
rect 766 812 829 924
rect 758 807 835 812
rect 758 406 768 807
rect 825 406 835 807
rect 758 401 835 406
rect 152 289 222 294
rect 841 289 917 292
rect 152 229 157 289
rect 217 287 917 289
rect 217 231 851 287
rect 907 231 917 287
rect 217 229 917 231
rect 152 224 222 229
rect 841 226 917 229
use sky130_fd_pr__pfet_01v8_2ZH9AN  sky130_fd_pr__pfet_01v8_2ZH9AN_0
timestamp 1729132718
transform 1 0 231 0 1 606
box -109 -262 109 262
use sky130_fd_pr__pfet_01v8_2ZH9AN  sky130_fd_pr__pfet_01v8_2ZH9AN_1
timestamp 1729132718
transform 1 0 231 0 1 -89
box -109 -262 109 262
use sky130_fd_pr__pfet_01v8_2ZH9AN  sky130_fd_pr__pfet_01v8_2ZH9AN_2
timestamp 1729132718
transform 1 0 835 0 1 -89
box -109 -262 109 262
use sky130_fd_pr__pfet_01v8_2ZH9AN  sky130_fd_pr__pfet_01v8_2ZH9AN_3
timestamp 1729132718
transform 1 0 835 0 1 606
box -109 -262 109 262
use sky130_fd_pr__pfet_01v8_2ZH9AN  sky130_fd_pr__pfet_01v8_2ZH9AN_4
timestamp 1729132718
transform 1 0 835 0 1 1301
box -109 -262 109 262
use sky130_fd_pr__pfet_01v8_2ZH9AN  sky130_fd_pr__pfet_01v8_2ZH9AN_5
timestamp 1729132718
transform 1 0 835 0 1 1996
box -109 -262 109 262
use sky130_fd_pr__pfet_01v8_2ZH9AN  sky130_fd_pr__pfet_01v8_2ZH9AN_6
timestamp 1729132718
transform 1 0 231 0 1 1996
box -109 -262 109 262
use sky130_fd_pr__pfet_01v8_2ZH9AN  sky130_fd_pr__pfet_01v8_2ZH9AN_7
timestamp 1729132718
transform 1 0 231 0 1 1301
box -109 -262 109 262
use sky130_fd_pr__pfet_01v8_SDE6B7  sky130_fd_pr__pfet_01v8_SDE6B7_0
timestamp 1729135886
transform 1 0 533 0 1 1996
box -323 -300 323 300
use sky130_fd_pr__pfet_01v8_SDE6B7  sky130_fd_pr__pfet_01v8_SDE6B7_1
timestamp 1729135886
transform 1 0 533 0 1 1301
box -323 -300 323 300
use sky130_fd_pr__pfet_01v8_SDE6B7  sky130_fd_pr__pfet_01v8_SDE6B7_2
timestamp 1729135886
transform 1 0 533 0 1 606
box -323 -300 323 300
use sky130_fd_pr__pfet_01v8_SDE6B7  sky130_fd_pr__pfet_01v8_SDE6B7_3
timestamp 1729135886
transform 1 0 533 0 1 -89
box -323 -300 323 300
<< labels >>
flabel metal3 782 862 782 862 0 FreeSans 800 0 0 0 D1
port 2 nsew
flabel metal1 878 2302 878 2302 0 FreeSans 800 0 0 0 VDD
port 4 nsew
flabel via1 792 1048 792 1048 0 FreeSans 800 0 0 0 D2
port 1 nsew
flabel metal2 880 904 880 904 0 FreeSans 800 0 0 0 D5
port 0 nsew
<< end >>
